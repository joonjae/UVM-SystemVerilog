interface uart_clk_if;
    logic clk, rst;
    logic [16:0] baund;
    logic tx_clk;
endinterface