module top (
  input [2:0] a, b,
  input rst,
  input feed,
  output [2:0] y,
  output done
);
  
/*
 
User Logic here
Do not add anything
..............
............
...........
.........
.......
 
*/
  
  endmodule